// Copyright Supranational LLC
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

`ifndef ADDER_DEFINES_SV
`define ADDER_DEFINES_SV

// Processors (white/gray/black)
localparam int W_P = 0;
localparam int G_P = 1;
localparam int B_P = 2;

`endif
